package common_pkg;
  parameter TEST_PARAM = 12;
  int test_int = 14;

  typedef struct packed {
    logic        a;
    logic        b;
  } mytype2_t;

endpackage // common_pkg
